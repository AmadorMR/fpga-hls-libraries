`timescale 1ns/100ps
module mipicsi2rxdecoderPF #(parameter g_DATAWIDTH = 10,
                             parameter g_LANE_WIDTH = 2,
                             parameter g_NUM_OF_PIXELS = 1,
                             parameter g_INPUT_DATA_INVERT = 0,
                             parameter g_BUFF_DEPTH = 1920)
                           (input CAM_CLOCK_I,
                            input PARALLEL_CLOCK_I,
                            input RESET_n_I,
                            input[7 : 0] L0_HS_DATA_I,
                            input[7 : 0] L1_HS_DATA_I,
                            input[7 : 0] L2_HS_DATA_I,
                            input[7 : 0] L3_HS_DATA_I,
                            input[7 : 0] L4_HS_DATA_I,
                            input[7 : 0] L5_HS_DATA_I,
                            input[7 : 0] L6_HS_DATA_I,
                            input[7 : 0] L7_HS_DATA_I,
                            input L0_LP_DATA_I,
                            input L0_LP_DATA_N_I,
                            input L1_LP_DATA_I,
                            input L1_LP_DATA_N_I,
                            input L2_LP_DATA_I,
                            input L2_LP_DATA_N_I,
                            input L3_LP_DATA_I,
                            input L3_LP_DATA_N_I,
                            input L4_LP_DATA_I,
                            input L4_LP_DATA_N_I,
                            input L5_LP_DATA_I,
                            input L5_LP_DATA_N_I,
                            input L6_LP_DATA_I,
                            input L6_LP_DATA_N_I,
                            input L7_LP_DATA_I,
                            input L7_LP_DATA_N_I,
                            output[g_NUM_OF_PIXELS * g_DATAWIDTH - 1 : 0] data_out_o,
                            output frame_end_o,
                            output frame_start_o,
                            output frame_valid_o,
                            output line_end_o,
                            output line_start_o,
                            output line_valid_o,
                            output[15 : 0] word_count_o);
  wire[7 : 0] lolI;
  wire[7 : 0] oolI;
  wire[7 : 0] iolI;
  wire[7 : 0] OilI;
  wire[7 : 0] IilI;
  wire[7 : 0] lilI;
  wire[7 : 0] oilI;
  wire[7 : 0] iilI;
  embsync_detect #(.g_LANE_WIDTH(g_LANE_WIDTH)) OO0I(.RESET_N_I(RESET_n_I),
                                                     .CLOCK_I(CAM_CLOCK_I),
                                                     .L0_DATA_I(L0_HS_DATA_I),
                                                     .L1_DATA_I(L1_HS_DATA_I),
                                                     .L2_DATA_I(L2_HS_DATA_I),
                                                     .L3_DATA_I(L3_HS_DATA_I),
                                                     .L4_DATA_I(L4_HS_DATA_I),
                                                     .L5_DATA_I(L5_HS_DATA_I),
                                                     .L6_DATA_I(L6_HS_DATA_I),
                                                     .L7_DATA_I(L7_HS_DATA_I),
                                                     .L0_LP_DATA_N_I(L0_LP_DATA_N_I),
                                                     .L1_LP_DATA_N_I(L1_LP_DATA_N_I),
                                                     .L2_LP_DATA_N_I(L2_LP_DATA_N_I),
                                                     .L3_LP_DATA_N_I(L3_LP_DATA_N_I),
                                                     .L4_LP_DATA_N_I(L4_LP_DATA_N_I),
                                                     .L5_LP_DATA_N_I(L5_LP_DATA_N_I),
                                                     .L6_LP_DATA_N_I(L6_LP_DATA_N_I),
                                                     .L7_LP_DATA_N_I(L7_LP_DATA_N_I),
                                                     .L0_DATA_O(lolI),
                                                     .L1_DATA_O(oolI),
                                                     .L2_DATA_O(iolI),
                                                     .L3_DATA_O(OilI),
                                                     .L4_DATA_O(IilI),
                                                     .L5_DATA_O(lilI),
                                                     .L6_DATA_O(oilI),
                                                     .L7_DATA_O(iilI));
  mipi_csi2_rxdecoder #(.g_DATAWIDTH(g_DATAWIDTH), .g_INPUT_DATA_INVERT(g_INPUT_DATA_INVERT), .g_LANE_WIDTH(g_LANE_WIDTH), .g_NUM_OF_PIXELS(g_NUM_OF_PIXELS), .g_BUFF_DEPTH(g_BUFF_DEPTH)) IO0I(.CAM_CLOCK_I(CAM_CLOCK_I),
                                                                                                                                                                                                .READ_CLOCK_I(PARALLEL_CLOCK_I),
                                                                                                                                                                                                .RESET_n_I(RESET_n_I),
                                                                                                                                                                                                .ChannelA_i(lolI),
                                                                                                                                                                                                .ChannelB_i(oolI),
                                                                                                                                                                                                .ChannelC_i(iolI),
                                                                                                                                                                                                .ChannelD_i(OilI),
                                                                                                                                                                                                .ChannelE_i(IilI),
                                                                                                                                                                                                .ChannelF_i(lilI),
                                                                                                                                                                                                .ChannelG_i(oilI),
                                                                                                                                                                                                .ChannelH_i(iilI),
                                                                                                                                                                                                .pixel_valid_o(line_valid_o),
                                                                                                                                                                                                .frame_start_o(frame_start_o),
                                                                                                                                                                                                .frame_end_o(frame_end_o),
                                                                                                                                                                                                .frame_valid_o(frame_valid_o),
                                                                                                                                                                                                .line_start_o(line_start_o),
                                                                                                                                                                                                .line_end_o(line_end_o),
                                                                                                                                                                                                .data_out_o(data_out_o),
                                                                                                                                                                                                .word_count_o(word_count_o),
                                                                                                                                                                                                .frame_number_o());
endmodule
